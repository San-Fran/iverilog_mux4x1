//mux4x1.v
//Author: Francisco Vega
//CSC 205

module MuxMod(s, s1, d0, d1, d2, d3, o);  // module definition
   input s, s1, d0, d1, d2, d3;
   output o;
  
   wire s_inv, s1_inv, and0, and1, and2, and3;
   
    not(s_inv, s);
    not(s1_inv, s1);
   
    and(and0, s_inv, s1_inv, d0);
    and(and1, s1_inv, s, d1);
    and(and2, s_inv, s1, d2);
    and(and3, s, s1, d3);
    or(o, and0, and1, and2, and3);
endmodule

module TestMod;   // module to test-run
   reg s, s1, d0, d1, d2, d3;       
   wire o;   

   MuxMod my_mux(s, s1, d0, d1, d2, d3, o); // create instance

   initial begin
      $monitor("%5d\t%b\t%b\t%b\t%b\t%b\t%b\t", $time, s1, s, d0, d1, d2, d3, o);
      $display(" Time\ts1\ts0\td0\td1\td2\td3\to");
      $display("-----------------------------------------------------------");
      #63;
      $finish;
   end

   always begin   // infinite loop
      s1 = 0; s = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;         // wait 1 simulation time unit/cycle
      s1 = 0; s = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 0; s = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0;
      #1;
      s1 = 1; s = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1;
      #1;
   end
endmodule

